module NpuExecuteController(
  input         clock,
  input         reset,
  output        io_cmd_ready, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input         io_cmd_valid, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input  [15:0] io_cmd_bits_aBase, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input  [15:0] io_cmd_bits_bBase, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input  [15:0] io_cmd_bits_cBase, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input         io_cmd_bits_start, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input         io_spR_0_req_ready, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output        io_spR_0_req_valid, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [7:0]  io_spR_0_req_bits, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input         io_spR_0_resp_valid, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input  [63:0] io_spR_0_resp_bits, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input         io_spR_1_req_ready, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output        io_spR_1_req_valid, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [7:0]  io_spR_1_req_bits, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input         io_spR_1_resp_valid, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input  [63:0] io_spR_1_resp_bits, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input         io_spR_2_req_ready, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output        io_spR_2_req_valid, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [7:0]  io_spR_2_req_bits, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input         io_spR_2_resp_valid, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input  [63:0] io_spR_2_resp_bits, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input         io_spR_3_req_ready, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output        io_spR_3_req_valid, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [7:0]  io_spR_3_req_bits, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input         io_spR_3_resp_valid, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input  [63:0] io_spR_3_resp_bits, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output        io_spW_0_en, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [7:0]  io_spW_0_addr, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [63:0] io_spW_0_data, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output        io_spW_1_en, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [7:0]  io_spW_1_addr, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [63:0] io_spW_1_data, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output        io_spW_2_en, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [7:0]  io_spW_2_addr, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [63:0] io_spW_2_data, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output        io_spW_3_en, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [7:0]  io_spW_3_addr, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [63:0] io_spW_3_data, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input         io_mesh_a_ready, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output        io_mesh_a_valid, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [63:0] io_mesh_a_bits, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input         io_mesh_b_ready, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output        io_mesh_b_valid, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output [63:0] io_mesh_b_bits, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input         io_mesh_d_valid, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  input  [63:0] io_mesh_d_bits, // @[src/main/scala/npu/ExecutionController.scala 52:14]
  output        io_done // @[src/main/scala/npu/ExecutionController.scala 52:14]
);


// Write your code here

endmodule
